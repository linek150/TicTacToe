library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

--AI PLAYER IS ALWAYS PLAYER CP='0'

--HUMAN PLAYER IS ON BOARD AS "11"


entity AI is
    Port (
    clk 	: in std_logic;
    rst 	: in std_logic;
    CP 		: in std_logic;--current player
	AIPAI	: in std_logic;--Artificial Intelligence player action iniciation
	AICB 	: in std_logic_vector(17 downto 0);
	AION	: in std_logic_vector(1 downto 0);
	AICL	: out std_logic_vector(8 downto 0);
	AIFCLR	:out std_logic
     );
end AI;

architecture Behav of AI is
type state is (waiting, move);
signal currentState:state;
type rotation is (one,two,three,four,five,six,none);
signal boardRotation	: rotation;
signal AIICL			: std_logic_vector(0 to 8);--AI internal Current LOcation 
signal AICLR			: std_logic_vector(8 downto 0);--AI internal Current LOcation 
signal IB 				:std_logic_vector(0 to 17);
signal CB 				:std_logic_vector(0 to 17);
signal AIFCLRIn         :std_logic;

begin
--downto and to change
CB<=AICB(0)&AICB(1)&AICB(2)&AICB(3)&AICB(4)&AICB(5)&AICB(6)&AICB(7)&AICB(8)&AICB(9)
	&AICB(10)&AICB(11)&AICB(12)&AICB(13)&AICB(14)&AICB(15)&AICB(16)&AICB(17);

--Board Rotation
process(clk,rst)
begin
	if rst='1' then
		boardRotation<=none;
	elsif rising_edge(clk) then
		if CB="000011000000000000" then
			boardRotation<=one;
		elsif CB="000000110000000000" then
			boardRotation<=two;
		elsif CB="000000000011000000" then 
			boardRotation<=three;
		elsif CB="000000000000110000" then
			boardRotation<=four;
		elsif CB="000000000000001100" then
			boardRotation<=five;
		elsif CB="000000000000000011" then 
			boardRotation<=six;
		elsif CB="000000000000000000" then		
			boardRotation<=none;
		end if;
	end if;
end process;
 
-- board rotation
IB<=CB when boardRotation=none else
	CB(4 to 5)&CB(2 to 3)&CB(0 to 1)&CB(10 to 11)&CB(8 to 9)&CB(6 to 7)&CB(16 to 17)&CB(14 to 15)&CB(12 to 13) when boardRotation=one else
	CB(0 to 1)&CB(6 to 7)&CB(12 to 13)&CB(2 to 3)&CB(8 to 9)&CB(14 to 15)&CB(4 to 5)&CB(10 to 11)&CB(16 to 17) when boardRotation=two else
	CB(4 to 5)&CB(10 to 11)&CB(16 to 17)&CB(2 to 3)&CB(8 to 9)&CB(14 to 15)&CB(0 to 1)&CB(6 to 7)&CB(12 to 13) when boardRotation=three else
	CB(12 to 17)&CB(6 to 11)&CB(0 to 5) when boardRotation=four else
	CB(12 to 17)&CB(6 to 11)&CB(0 to 5)	when boardRotation=five else 
	CB(16 to 17)&CB(10 to 11)&CB(4 to 5)&CB(14 to 15)&CB(8 to 9)&CB(2 to 3)&CB(12 to 13)&CB(6 to 7)&CB(0 to 1) when boardRotation=six else
	(others=>'0');
	
--AIICL rotation based on current rotation state
AICLR<=AIICL when boardRotation=none else
	AIICL(2)&AIICL(1)&AIICL(0)&AIICL(5)&AIICL(4)&AIICL(3)&AIICL(8)&AIICL(7)&AIICL(6)  when boardRotation=one else	
	AIICL(0)&AIICL(3)&AIICL(6)&AIICL(1)&AIICL(4)&AIICL(7)&AIICL(2)&AIICL(5)&AIICL(8) when boardRotation=two else
	AIICL(6)&AIICL(3)&AIICL(0)&AIICL(7)&AIICL(4)&AIICL(1)&AIICL(8)&AIICL(5)&AIICL(2) when boardRotation=three else
	AIICL(6)&AIICL(7)&AIICL(8)&AIICL(3)&AIICL(4)&AIICL(5)&AIICL(0)&AIICL(1)&AIICL(2) when boardRotation =four or boardRotation=five else
	AIICL(8)&AIICL(5)&AIICL(2)&AIICL(7)&AIICL(4)&AIICL(1)&AIICL(6)&AIICL(3)&AIICL(0) when boardRotation=six else
	(others=>'0');

AICL<=AICLR(0)&AICLR(1)&AICLR(2)&AICLR(3)&AICLR(4)&AICLR(5)&AICLR(6)&AICLR(7)&AICLR(8);
	
	
	
--100000000000000000
--AI move based on Current Board
process(clk,rst)
begin

	if rst='1' then
		AIICL<=(others=>'0');
	elsif rising_edge(clk) then
		if AIPAI='1' and CP='0' and AION="11" then
			if  
			IB="001111001000000000" or IB="001100111000000000" or IB="001100001000001100" or IB="001111101011110010" or
			IB="001100101011111110" or IB="001110001011110000" or IB="001111111010100011" or IB="000000001100000000" or 
			IB="000000000000000000"
			then --0
				AIICL<="100000000";
                
				
			elsif
			IB="110011001000000000"	or IB="110011111000100000" or IB="110000101011110000" or IB="110011111010101100" or
			IB="100000001100001100" or IB="100011111110101100" or IB="100011111110100011" or IB="100000111110001100" or 
			IB="100010111110110011" or IB="100010111110001111" or IB="100010101111111100" or IB="100010101111110011" or 
			IB="100010111100110000" or IB="100010001111110000" or IB="100010001100111100" or IB="100010001100110011" or --16
			IB="100000111110101111" or IB="100011111010111011" or IB="100011111010101111" or IB="100010101111110000" or --20
			IB="100010101100111100" or IB="100010101100110011" or IB="100010001011110011" or IB="100011001000111011" or 
			IB="100000111000111011" or IB="100000001011111011" or IB="100010110000000011" or IB="100010001100000011" or	--28
			IB="100010000011000011" or IB="100010000000110011" or IB="100010000000001111"
			then--1 
				AIICL<="010000000";
                
				
			elsif
			IB="111100001000000000" or IB="110000001011000000" or IB="111100111000100000" or IB="110000111011100000" or
			IB="110000111000101100" or IB="110000111000100011" or IB="111100111010101100" or IB="110000111010101111" or 
			IB="110000101011000011" or IB="111100001000000000" or IB="001100001011000000" or IB="101100111011100011" or
			IB="101100111000101111" or IB="111100101011110010" or IB="101100001011101111" or IB="111100111010100011" or 
			IB="001100111010101111" or IB="100000001100110000" or IB="101100001100111000" or IB="101100111110111000" or --20
			IB="101100101111111000" or IB="101100101100111011" or IB="100000111110110000" or IB="100000111110000011" or
			IB="101000111110111100" or IB="101000111110001111" or IB="100000101111110000" or IB="101000111100001100" or --28
			IB="101000001111001100" or IB="101000001100111100" or IB="101000001100001111" or IB="100000000000000011" or --32
			IB="101100001000000011" or IB="101100111000100011" or IB="100000111011100011" or IB="100000111000101111" or --36
			IB="100000101100110000" or IB="100000001011000011" or IB="101100111010111011" or IB="101100001000101111" or --40
			IB="100000001011101111"
			then--2
				AIICL<="001000000";
                
				
			elsif 
			IB="110000001000110000" or IB="110000001000000011" or IB="111110001000110000" or IB="110010001011110000" or
			IB="111100001010001100" or IB="110011001010001100" or IB="110000001010111100" or IB="110000001010001111" or
			IB="001100001000110000" or IB="111110001000110000" or IB="111100001010000011" or IB="001111001010000011" or 
			IB="001100001010110011" or IB="001100001010001111" or IB="100000001111000000" or IB="101100001111001000" or 
			IB="101100001100001011" or IB="101111001100101011" or IB="101110001111111000" or IB="101110001100111011" or
			IB="101111001100100000" or IB="100011001111100000" or IB="100011001100101100" or IB="100011001100100011" or	--24
			IB="101011001111101100" or IB="101011001100101111" or IB="101100001100100011" or IB="100000001111100011" or --28
			IB="100000001100101111" or IB="100000001100000000" or IB="101110001011111011" or IB="101111001010000011" or 
			IB="100011001010110011" or IB="100011001010001111" or IB="101111001010111011" or IB="100011001000101111" or	--36
			IB="101110001100100011" or IB="101110000011100011" or IB="101110000000101111"
			then--3
				AIICL<="000100000";
                
				
			elsif
			IB="110000000000000000" or IB="001100000000000000" or IB="101100000000000000" or IB="100011000000000000" or 
			IB="100000110000000000" or IB="100000000011000000" or IB="100000000000110000" or IB="100000000000001100" or 
			IB="101110110000100011" 
			then--4
				AIICL<="000010000";
                
				
			elsif 
			IB="110000001000001100" or IB="111110101000111100" or IB="111110101000110011" or IB="111011111000101100" or
			IB="111011001000101111" or IB="111011111000101100" or IB="111100101000110000" or IB="110011101000110000" or 
			IB="110000101000111100" or IB="110000101000110011" or IB="111100101000000011" or IB="110011101000000011" or 
			IB="110000101000110011" or IB="110000101000001111" or IB="001100001000000011" or IB="111110101000111100" or
			IB="111110101000110011" or IB="101111001000000011" or IB="101111111000100011" or IB="111100111000110000" or
			IB="001111101000110000" or IB="001100101000111100" or IB="001100101000110011" or IB="101111001000101111" or--24
			IB="100000111100000000" or IB="101100111100001000" or IB="101110111100111000" or IB="100011111100100000" or--28
			IB="101011111100101100" or IB="100000111100100011" or IB="101110111000111011" or IB="100011001000000011" or--32
			IB="100011111000100011" or IB="101110101100111011" or IB="101100001000111011"
			then--5
				AIICL<="000001000";
                
				
			elsif 
			IB="110000111000000000" or IB="001110111000000000" or IB="111110001011000000" or IB="111110001000001100" or 
			IB="111110001000000011" or IB="111011001000001100" or IB="111110001011000000" or IB="110010111011000000" or
			IB="110010001011001100" or IB="110010001011000011" or IB="110000111010001100" or IB="111110101011000011" or 
			IB="110010101011001111" or IB="111110111000000000" or IB="111110001011000000" or IB="111110001000001100" or
			IB="111110001000000011" or IB="101100111000000011" or IB="111110001011000000" or IB="001110111011000000" or 
			IB="001110001011001100" or IB="001110001011000011" or IB="101100001000001111" or IB="001100111010000011" or --24
			IB="100011001100000000" or IB="100000001100000011" or IB="101111001100001000" or IB="101111111110001000" or 
			IB="101100111110001011" or IB="101111101111001000" or IB="101100101111001011" or IB="101111101100001011" or	--32
			IB="100011111110000000" or IB="101011111110001100" or IB="101100101111000000" or IB="100011101111000000" or --36
			IB="100000101111001100" or IB="100000101111000011" or IB="101011001100001100" or IB="101110111000000011" or --40
			IB="101110001011000011" or IB="101110001000001111" or IB="101111111010001011" or IB="100000111000000011" or	--44
			IB="101100101100000000" or IB="100011101100000000" or IB="100000101111000000" or IB="100000101100001100" or --48
			IB="100000101100000011" or IB="100010111011000011" or IB="100010001011001111" or IB="100000001000001111" or --52
			IB="101110000000000011"
			then--6
				AIICL<="000000100";
                
				
			elsif
			IB="111110101011110000" or IB="111011111000000000" or IB="111011001011000000" or IB="111011001000110000" or
			IB="111011001000000011" or IB="111011111011100000" or IB="111011111000100011" or IB="111110101011110000" or
			IB="110010101011110011" or IB="111011101011110000" or IB="111000101011110011" or IB="110010101011110011" or
			IB="111110101011110000" or IB="101110001011110011" or IB="101100001100000000" or IB="101111111110100000" or 
			IB="101100111110000000" or IB="101110111110000011" or IB="101110101111110000" or IB="101110001100110000" or	--20
			IB="101100111110100011" or IB="101110001000110011" or IB="100011111010000011" or IB="101111111010100011" or	--24
			IB="101110101100110000" or IB="100000001000110011"
			then--7
				AIICL<="000000010";
			    
			
			elsif
			IB="111011001011101100" or IB="110010101011111100" or IB="111000101011111100" or IB="101111111000000000" or
			IB="101111001011000000" or IB="101111001000110000" or IB="101111001000001100" or IB="101111111000000000" or
			IB="101100111011000000" or IB="101100111000110000" or IB="101100111000001100" or IB="001100101011110000" or 
			IB="101110111011110000" or IB="101110001011111100" or IB="101100001011001100" or IB="101100001000111100" or 
			IB="101111111100101000" or IB="101111001111101000" or IB="101110111110110000" or IB="100010111110111100" or	--20
			IB="101111001000000000" or IB="101100111000000000" or IB="101100001011000000" or IB="101100001000110000" or	--24
			IB="101100001000001100" or IB="100011111000000000" or IB="100011001011000000" or IB="100011001000110000" or	--28
			IB="100011001000001100" or IB="100000111011000000" or IB="100000111000110000" or IB="100000111000001100" or --32
			IB="101110101111111000" or IB="100000001011110000" or IB="100000001011001100" or IB="100000001000111100" 	--36
			then--8
				AIICL<="000000001";
				
			end if;	
			AIFCLR<='1';
		else
			AIFCLR<='0';
			AIICL<=(others=>'0');
			end if;
	end if;
end process;
			
				
	
   
end Behav;
